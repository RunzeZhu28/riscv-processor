module control(

);

endmodule