module execution(

);
endmodule