module control(

);

endmodule
